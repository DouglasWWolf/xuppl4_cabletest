
//================================================================================================
//    Date      Vers   Who  Changes
// -----------------------------------------------------------------------------------------------
// 06-Dec-2023  1.0.0  DWW  Initial creation
//
// 05-May-2024  1.1.0  DWW  Added revision tracking
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 1;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;

localparam VERSION_DAY   = 5;
localparam VERSION_MONTH = 5;
localparam VERSION_YEAR  = 2024;

localparam RTL_TYPE      = 741776;
localparam RTL_SUBTYPE   = 0;
