/*
================================================================================================
  Vers     Date    Who  Changes
------- ----------------------------------------------------------------------------------------
 1.0.0  06-Dec-23  DWW  Initial creation
                                 
 1.1.0  05-May-24  DWW  Added revision tracking
                                      
 1.2.0  28-May-24  DWW  Updated to latest cmac_control in order to be able to configure
                        pre-emphasis on the CMAC serdes.
                                       
 1.3.0  08-Jun-24  DWW  Added run-time control over RS-FEC and the pre-emphasis setting
                                  
 1.4.0  15-Jun-24  DWW  Now controlling CMAC gt_txdiffctrl
                                    
 1.5.0  16-Jun-24  DWW  Added programmable gt_txpostcursor and gt_txdiffctrl
                                 
 1.5.1  30-Jun-24  DWW  Set SYSTEM_JITTER to 300ps to tighten up timing
                                  
 1.6.0  29-Nov-24  DWW  Added ILAs on the CMAC tx and rx streams
                                           
 1.8.0  04-Jul-25  DWW  Integrated with the build system
================================================================================================
*/

localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 8;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;


localparam RTL_TYPE      = 741776;
localparam RTL_SUBTYPE   = 0;
